library verilog;
use verilog.vl_types.all;
entity check_edge_tb is
end check_edge_tb;
