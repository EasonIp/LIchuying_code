library verilog;
use verilog.vl_types.all;
entity pll_tb is
end pll_tb;
