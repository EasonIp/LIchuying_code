`timescale 1ns/1ps

module adder_half_tb;

	reg a, b;
	
	wire sum;
	wire c_out;



endmodule
