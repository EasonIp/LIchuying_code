library verilog;
use verilog.vl_types.all;
entity iic_noack_tb is
end iic_noack_tb;
