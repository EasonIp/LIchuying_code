library verilog;
use verilog.vl_types.all;
entity ledrun_tb is
    generic(
        T1s             : integer := 5
    );
end ledrun_tb;
