library verilog;
use verilog.vl_types.all;
entity ledrun_tb is
end ledrun_tb;
