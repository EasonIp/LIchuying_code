library verilog;
use verilog.vl_types.all;
entity key_pad_tb is
end key_pad_tb;
