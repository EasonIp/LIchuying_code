library verilog;
use verilog.vl_types.all;
entity ps2_tb is
end ps2_tb;
