library verilog;
use verilog.vl_types.all;
entity divider2_tb is
end divider2_tb;
