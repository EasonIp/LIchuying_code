library verilog;
use verilog.vl_types.all;
entity seg7_tb is
end seg7_tb;
