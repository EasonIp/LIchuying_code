`timescale 1ns/1ps

module divider2_tb;

	reg clk, rst_n;
	
	wire clk_out;

	divider2 #(.WIDTH(6)) dut (.clk(clk), .rst_n(rst_n), .clk_out(clk_out));

	initial
		begin
			clk = 1;
			rst_n = 0;
			#200.1
			rst_n = 1;
			
			#500 $stop;
		end

	always #10 clk = ~clk;

endmodule
