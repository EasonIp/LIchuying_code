library verilog;
use verilog.vl_types.all;
entity adc_tb is
end adc_tb;
