library verilog;
use verilog.vl_types.all;
entity vga_tb is
end vga_tb;
