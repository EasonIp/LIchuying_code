library verilog;
use verilog.vl_types.all;
entity key_flag_tb is
end key_flag_tb;
