module top (clk, rst_n, key, r, g, b, hsync, vsync, VGA_CLK, VGA_BLANK, VGA_SYNC);

	input clk, rst_n;
	input [1:0] key;
	
	output [9:0] r, g, b;
	output hsync, vsync;
	output VGA_CLK;
	output VGA_BLANK, VGA_SYNC;
	
	assign VGA_BLANK = 1'b1;
	assign VGA_SYNC = 1'b0;
	
	wire [1:0] key_out;
	wire [29:0] rgb30;	
	wire [7:0] addr;
	wire [7:0] sine_q, square_q;
	wire [7:0] o_wave;

	parameter T20ms = 800_000;
	
	pll pll (.areset(~rst_n), .inclk0(clk), .c0(VGA_CLK));		// VGA_CLK is 40M clock

	jitter_key #(.T20ms(T20ms)) k1(
			.clk(VGA_CLK),
			.rst_n(rst_n),
			.key(key[0]), 
			.key_out(key_out[0])
		);  

	jitter_key #(.T20ms(T20ms)) k2(
			.clk(VGA_CLK),
			.rst_n(rst_n),
			.key(key[1]), 
			.key_out(key_out[1])
		);  
	
	sine_rom256	sine_rom256_inst (
			.address ( addr ),
			.clock ( VGA_CLK ),
			.q ( sine_q )
		);

	square_rom256	square_rom256_inst (
			.address ( addr ),
			.clock ( VGA_CLK ),
			.q ( square_q )
		);

	dds_controller ctrl(
			.clk(VGA_CLK), 
			.rst_n(rst_n), 
			.key_out(key_out), 
			.addr(addr), 
			.sine_q(sine_q), 
			.square_q(square_q), 
			.o_wave(o_wave)
		);

	vga_dds vga_dds (
			.clk(VGA_CLK), 
			.rst_n(rst_n), 
			.key_out(key_out), 
			.wave(o_wave), 
			.rgb30(rgb30), 
			.hsync(hsync), 
			.vsync(vsync)
		);
	
	rgb rgb (.rgb30(rgb30), .r(r), .g(g), .b(b));

endmodule
