library verilog;
use verilog.vl_types.all;
entity rca_16_tb is
end rca_16_tb;
